library verilog;
use verilog.vl_types.all;
entity tb_fpmul is
end tb_fpmul;
